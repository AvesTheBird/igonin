library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity adder is
  port (
    X1 : in std_logic
  );
end adder;

architecture rtl of circuit is
  signal and_2 : std_logic;
  signal not_6 : std_logic;
begin
end rtl;